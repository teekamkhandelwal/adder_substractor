interface simple (input logic clk, reset);
  logic load;
  logic load1;
  logic [3:0] a;
  logic [3:0] b;
  logic [4:0] sum;
  logic [4:0] sub;
  
endinterface
